`ifndef MONITOR_SVH
`define MONITOR_SVH
`include "uvm_macros.svh"
import uvm_pkg::*;

class common_cfg extends uvm_object;
        
endclass