package package_;
    `include "transaction.sv"
    `include "sequence.sv"
    `include "sequencer.sv"
    `include "driver.sv"
    `include "monitor.sv"
    `include "scoreboard.sv"
    `include "coverage.sv"
    `include "agent.sv"
    `include "env.sv"
    `include "test.sv"
    `include "common_cfg.sv"
endpackage