interface intf;
  logic         clk;
  logic         rst_n;
  logic  [7:0]  data_in0;
  logic  [7:0]  data_in1;
  logic  [7:0]  data_in2;
  logic  [7:0]  data_in3;
  logic         valid_in0;
  logic         valid_in1;
  logic         valid_in2;
  logic         valid_in3;
  logic  [7:0]  data_out0;
  logic  [7:0]  data_out1;
  logic         valid_out0;
  logic         valid_out1;
endinterface
